module top (
    input wire clk,
    input wire reset,
    input wire rx,
    output wire tx,
    output wire [5:0] led,
    inout [4:0]gpios
);



endmodule
