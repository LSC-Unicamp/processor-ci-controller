module top (
    input wire clk, // 50mhz clock
    output wire led
);


    
endmodule