module Interpreter #(
    parameter CLK_FREQ = 25000000
) (
    input wire clk,
    input wire reset
);
    
endmodule
